../../eth_test/src/udp_wrapper.vhd